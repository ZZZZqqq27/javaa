//IF/ID
//32+32+32
/*
module IFIDRegister(input clk,reset,clear,
input []

    )
    endmodule*/
//ID/EX
//20+32+32+32 +5+32+32
//第三第四间长度
//
//第四第五间长度

/*module floprc #(parameter WIDTH = 8)
              (input                  clk, reset, clear,
               input      [WIDTH-1:0] d, 
               output reg [WIDTH-1:0] q);

  always @(posedge clk, posedge reset)
    if (reset)      q <= 0;
    else if (clear) q <= 0;
    else            q <= d;
endmodule*/







